// Main state coding
parameter INIT_STATE            = 3'd0;
parameter ONLED0_15_STATE       = 3'd1;
parameter OFFLED15_5_STATE      = 3'd2;
parameter ONLED5_10_STATE       = 3'd3;
parameter OFFLED10_0_STATE      = 3'd4;
parameter ONLED0_5_STATE        = 3'd5;
parameter OFFLED5_0_STATE       = 3'd6;

// Counting encode
parameter COUNT_DIS             = 2'd0;
parameter COUNT_UP_EN           = 2'd1;
parameter COUNT_DOWN_EN         = 2'd2;

// Counter init value
parameter COUNTER_INIT          = 5'd0;

